module adder_div(dataa, datab, sum);

input [15:0] dataa; 
input datab;
output [15:0] sum; 

assign sum = dataa + datab;

endmodule 